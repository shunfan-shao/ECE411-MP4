package cpu_types;

// typedef struct packed {
//     rv32i_opcode opcode;
//     alu_ops aluop;
//     logic regfilemux_sel;
//     logic load_regfile;
//     /* ... other signals ... */
// } rv32i_control_word;



endpackage : cpu_types